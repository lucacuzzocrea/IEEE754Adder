library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ShiftRight48 is
	
	port(
		N : in std_logic_vector(47 downto 0);
		PLACES : in std_logic_vector(8 downto 0);
		RESULT : out std_logic_vector(47 downto 0)
	);

end ShiftRight48;


architecture ShiftRightArch of ShiftRight48 is

begin

	asdf: process (N, PLACES)
	
	begin
	
		case PLACES is
			when "000000000" => RESULT <= N( 47 downto 0 );
			when "000000001" => RESULT <= "0" & N( 47 downto 1 );
			when "000000010" => RESULT <= "00" & N( 47 downto 2 );
			when "000000011" => RESULT <= "000" & N( 47 downto 3 );
			when "000000100" => RESULT <= "0000" & N( 47 downto 4 );
			when "000000101" => RESULT <= "00000" & N( 47 downto 5 );
			when "000000110" => RESULT <= "000000" & N( 47 downto 6 );
			when "000000111" => RESULT <= "0000000" & N( 47 downto 7 );
			when "000001000" => RESULT <= "00000000" & N( 47 downto 8 );
			when "000001001" => RESULT <= "000000000" & N( 47 downto 9 );
			when "000001010" => RESULT <= "0000000000" & N( 47 downto 10 );
			when "000001011" => RESULT <= "00000000000" & N( 47 downto 11 );
			when "000001100" => RESULT <= "000000000000" & N( 47 downto 12 );
			when "000001101" => RESULT <= "0000000000000" & N( 47 downto 13 );
			when "000001110" => RESULT <= "00000000000000" & N( 47 downto 14 );
			when "000001111" => RESULT <= "000000000000000" & N( 47 downto 15 );
			when "000010000" => RESULT <= "0000000000000000" & N( 47 downto 16 );
			when "000010001" => RESULT <= "00000000000000000" & N( 47 downto 17 );
			when "000010010" => RESULT <= "000000000000000000" & N( 47 downto 18 );
			when "000010011" => RESULT <= "0000000000000000000" & N( 47 downto 19 );
			when "000010100" => RESULT <= "00000000000000000000" & N( 47 downto 20 );
			when "000010101" => RESULT <= "000000000000000000000" & N( 47 downto 21 );
			when "000010110" => RESULT <= "0000000000000000000000" & N( 47 downto 22 );
			when "000010111" => RESULT <= "00000000000000000000000" & N( 47 downto 23 );
			when "000011000" => RESULT <= "000000000000000000000000" & N( 47 downto 24 );
			when "000011001" => RESULT <= "0000000000000000000000000" & N( 47 downto 25 );
			when "000011010" => RESULT <= "00000000000000000000000000" & N( 47 downto 26 );
			when "000011011" => RESULT <= "000000000000000000000000000" & N( 47 downto 27 );
			when "000011100" => RESULT <= "0000000000000000000000000000" & N( 47 downto 28 );
			when "000011101" => RESULT <= "00000000000000000000000000000" & N( 47 downto 29 );
			when "000011110" => RESULT <= "000000000000000000000000000000" & N( 47 downto 30 );
			when "000011111" => RESULT <= "0000000000000000000000000000000" & N( 47 downto 31 );
			when "000100000" => RESULT <= "00000000000000000000000000000000" & N( 47 downto 32 );
			when "000100001" => RESULT <= "000000000000000000000000000000000" & N( 47 downto 33 );
			when "000100010" => RESULT <= "0000000000000000000000000000000000" & N( 47 downto 34 );
			when "000100011" => RESULT <= "00000000000000000000000000000000000" & N( 47 downto 35 );
			when "000100100" => RESULT <= "000000000000000000000000000000000000" & N( 47 downto 36 );
			when "000100101" => RESULT <= "0000000000000000000000000000000000000" & N( 47 downto 37 );
			when "000100110" => RESULT <= "00000000000000000000000000000000000000" & N( 47 downto 38 );
			when "000100111" => RESULT <= "000000000000000000000000000000000000000" & N( 47 downto 39 );
			when "000101000" => RESULT <= "0000000000000000000000000000000000000000" & N( 47 downto 40 );
			when "000101001" => RESULT <= "00000000000000000000000000000000000000000" & N( 47 downto 41 );
			when "000101010" => RESULT <= "000000000000000000000000000000000000000000" & N( 47 downto 42 );
			when "000101011" => RESULT <= "0000000000000000000000000000000000000000000" & N( 47 downto 43 );
			when "000101100" => RESULT <= "00000000000000000000000000000000000000000000" & N( 47 downto 44 );
			when "000101101" => RESULT <= "000000000000000000000000000000000000000000000" & N( 47 downto 45 );
			when "000101110" => RESULT <= "0000000000000000000000000000000000000000000000" & N( 47 downto 46 );
			when "000101111" => RESULT <= "00000000000000000000000000000000000000000000000" & N( 47 );
			when others   => RESULT <= "000000000000000000000000000000000000000000000000";
		end case;
		
	end process;

end ShiftRightArch;
